module single_port_ram(
    input data,
    input addr,
    input clk,
    input reset,
    output wdata
);

