module tb_piso_register();
    reg  clk,
    reg reset,
    reg load,
    reg [3:0] d,
    wire q


endmodule