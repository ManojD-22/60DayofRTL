module serial_in_parallel_out(
    input 
    );
endmodule