module piso_register(

    input clk,
    input reset,
    input [3:0] d,
    output reg q
);

endmodule